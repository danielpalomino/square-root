LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY square_root IS
	GENERIC (n: INTEGER:=8);
	PORT(
		clk, reset, start:	IN STD_LOGIC;
		number:		IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		pronto:			OUT STD_LOGIC;
		root:			OUT STD_LOGIC_VECTOR((n-1)/2 DOWNTO 0)
	);

END square_root;

ARCHITECTURE behavioral OF square_root IS

COMPONENT po  IS
	GENERIC (n: INTEGER:=8);
	PORT(
		clk, reset, start: IN STD_LOGIC;
		en_r, en_s, en_d, en_t, en_s_neg, en_clk: IN STD_LOGIC;
		number: IN STD_LOGIC_VECTOR (n-1 DOWNTO 0);
		mux0, mux1: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		mux_s: IN STD_LOGIC;
		ready: OUT STD_LOGIC;
		root: OUT STD_LOGIC_VECTOR (n-1 DOWNTO 0)
	);

END COMPONENT;

COMPONENT pc IS
	PORT(
		clk, reset, ready, start: IN STD_LOGIC;
		start_po, en_r, en_s, en_d, en_t, en_s_neg, en_clk, pronto: OUT STD_LOGIC;
		mux0, mux1: OUT STD_LOGIC_VECTOR (1 DOWNTO 0 );
		mux_s: OUT STD_LOGIC
	);

END COMPONENT;

SIGNAL reg_number, temp_root: STD_LOGIC_VECTOR (n-1 DOWNTO 0);
SIGNAL start_po, en_r, en_s, en_d, en_t, en_s_neg, en_clk, ready: STD_LOGIC;
SIGNAL mux0, mux1: STD_LOGIC_VECTOR (1 DOWNTO 0 );
SIGNAL mux_s: STD_LOGIC;

BEGIN

PROCESS (clk, reset)
BEGIN
	IF reset = '1' THEN
		reg_number <= (OTHERS=>'0');
		root <= (OTHERS=>'0');
	ELSIF clk'EVENT AND clk='1' THEN
		reg_number <= number;
		root <= temp_root((n-1)/2 DOWNTO 0);
	END IF;
END PROCESS;

PARTE_OPERATIVA: po GENERIC MAP (n) PORT MAP (
clk => clk,
reset => reset,
start => start_po,
en_r => en_r,
en_s => en_s,
en_d => en_d,
en_t => en_t,
en_s_neg => en_s_neg,
en_clk => en_clk,
number => reg_number,
mux0 => mux0,
mux1 => mux1,
mux_s => mux_s,
ready => ready,
root => temp_root
);

PARTE_CONTROLE: pc PORT MAP (
clk => clk,
reset => reset,
ready => ready,
start => start,
start_po => start_po,
en_r => en_r,
en_s => en_s,
en_d => en_d,
en_t => en_t,
en_s_neg => en_s_neg,
en_clk => en_clk,
pronto => pronto,
mux0 => mux0,
mux1 => mux1,
mux_s => mux_s
);
	
END behavioral;